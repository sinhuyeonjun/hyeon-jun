module tlqkf(
    in_a,
    out
);

input [2:0] in_a;
output reg [2:0]out;


endmodule 
library verilog;
use verilog.vl_types.all;
entity multiplexer is
    port(
        in_0            : in     vl_logic;
        in_1            : in     vl_logic;
        in_2            : in     vl_logic;
        in_3            : in     vl_logic;
        inx_4           : in     vl_logic;
        inx_5           : in     vl_logic;
        \out\           : out    vl_logic
    );
end multiplexer;

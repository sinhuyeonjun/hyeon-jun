library verilog;
use verilog.vl_types.all;
entity encoder is
    port(
        in_0            : in     vl_logic;
        in_1            : in     vl_logic;
        in_2            : in     vl_logic;
        in_3            : in     vl_logic;
        in_4            : in     vl_logic;
        in_5            : in     vl_logic;
        in_6            : in     vl_logic;
        in_7            : in     vl_logic;
        out_a           : out    vl_logic;
        out_b           : out    vl_logic;
        out_c           : out    vl_logic
    );
end encoder;
